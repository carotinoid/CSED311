module PC(
    input reset,
    input clk,
    input [31:0] next_pc,
    output [31:0] current_pc
);

endmodule