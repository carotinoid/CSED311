`include "vending_machine_def.v"

module calc_total(current_total, i_input_coin, coin_value, next_total);

    input current_total;
    input [`kNumCoins-1:0] i_input_coin;
    input 

    always @(*) begin
        next_total = current_total;
    
    end

endmodule